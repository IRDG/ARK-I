------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BasicPackage.ALL;
USE WORK.AluPackage  .ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY PartialProduct IS
    
    PORT   (A  : IN  uint32;
            B  : IN  uint32;
            PP : OUT PartialProductT
           );

END ENTITY PartialProduct;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE MainArch OF PartialProduct IS

SIGNAL SpecB : PartialProductT;

BEGIN

----------------------------------------------------------
-- 
-- Calculate partial products using AND gates
-- 
----------------------------------------------------------

IterateB: FOR I IN 0 TO 31 GENERATE
    
    SpecB(I) <= (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I)) &
                (B(I));
    
    PP(I) <= A AND SpecB(I);
    
END GENERATE IterateB;

END MainArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.PartialProduct(MainArch)
--PORT MAP   (A  => SLV,
--            B  => SLV,
--            PP => SLV
--           );
------------------------------------------------------------------------------------------