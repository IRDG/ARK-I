------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

USE WORK.BasicPackage.ALL;

ENTITY S1DecodeStageTestProtocol IS
END S1DecodeStageTestProtocol;

ARCHITECTURE S1DecodeStageTestProtocolArch OF S1DecodeStageTestProtocol IS

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------



BEGIN



END S1DecodeStageTestProtocolArch;
