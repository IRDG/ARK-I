------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BasicPackage.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY LocalClockModule IS
    
    PORT   (ClkConfig : IN  STD_LOGIC;
            Rst       : IN  STD_LOGIC;
            Clk       : IN  STD_LOGIC;
            LocalClk  : OUT STD_LOGIC
           );
    
END ENTITY LocalClockModule;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE MainArch OF LocalClockModule IS

BEGIN

------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------

LocalClk <= Clk;

END MainArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.LocalClockModule(MainArch)
--PORT MAP   (ClkConfig => SLV,
--            Rst       => SLV,
--            Clk       => SLV,
--            LocalClk  => SLV
--           );
------------------------------------------------------------------------------------------