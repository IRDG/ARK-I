------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY FullAdderHalfAdder IS
    
    PORT   (A    : IN  STD_LOGIC;
            B    : IN  STD_LOGIC;
            Cin  : IN  STD_LOGIC;
            R    : OUT STD_LOGIC;
            Cout : OUT STD_LOGIC
           );

END ENTITY FullAdderHalfAdder;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE FullAdder OF FullAdderHalfAdder IS

SIGNAL Mid : STD_LOGIC;

BEGIN

Mid  <=  A   XOR B  ;
R    <=  Mid XOR Cin;
Cout <= (A   AND B  ) OR (Mid AND Cin);

END FullAdder;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE HalfAdder OF FullAdderHalfAdder IS

BEGIN

R    <= A XOR B;
Cout <= A AND B;

END HalfAdder;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.FullAdderHalfAdder(FullAdder HalfAdder)
--PORT MAP   (A    => SLV,
--            B    => SLV,
--            Cin  => SLV,
--            R    => SLV,
--            Cout => SLV
--           );
------------------------------------------------------------------------------------------