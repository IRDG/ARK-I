------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

USE WORK.BasicPackage.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY Comparator IS
    
    PORT   (A           : IN  uint32;
            B           : IN  uint32;
            Comparisson : OUT uint06 
           );
    
END ENTITY Comparator;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE MainArch OF Comparator IS

BEGIN

------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------

Comparisson(0) <= '1' WHEN  (  SIGNED(A)  >   SIGNED(B))                                 ELSE
                  '0';

Comparisson(1) <= '1' WHEN  (  SIGNED(A)  <   SIGNED(B))                                 ELSE
                  '0';

Comparisson(2) <= '1' WHEN  (UNSIGNED(A)  = UNSIGNED(B))                                 ELSE
                  '0';

Comparisson(3) <= '1' WHEN ((UNSIGNED(A)  > UNSIGNED(B)) OR (UNSIGNED(A) < UNSIGNED(B))) ELSE
                  '0';

Comparisson(4) <= '1' WHEN  (UNSIGNED(A)  > UNSIGNED(B))                                 ELSE
                  '0';

Comparisson(5) <= '1' WHEN  (UNSIGNED(A)  < UNSIGNED(B))                                 ELSE
                  '0';

END MainArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.Comparator(MainArch)
--PORT MAP   (A           => SLV,
--            B           => SLV,
--            Comparisson => SLV
--           );
------------------------------------------------------------------------------------------