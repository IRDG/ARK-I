------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BasicPackage.ALL;
USE WORK.CachePackage.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY CacheOutputDecoder IS
    
    PORT   (Miss         : IN  SliceVectorT;
            RdDataArray  : IN  RdDataArrayT;
            SliceDataOut : OUT uint32       
           );
    
END ENTITY CacheOutputDecoder;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE MainArch OF CacheOutputDecoder IS

SIGNAL DecodedMiss : STD_LOGIC_VECTOR(SliceSize-1 DOWNTO 0);

BEGIN

------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------

WITH Miss SELECT
DecodedMiss <= x"0" WHEN "1111111111111110",
               x"1" WHEN "1111111111111101",
               x"2" WHEN "1111111111111011",
               x"3" WHEN "1111111111110111",
               x"4" WHEN "1111111111101111",
               x"5" WHEN "1111111111011111",
               x"6" WHEN "1111111110111111",
               x"7" WHEN "1111111101111111",
               x"8" WHEN "1111111011111111",
               x"9" WHEN "1111110111111111",
               x"A" WHEN "1111101111111111",
               x"B" WHEN "1111011111111111",
               x"C" WHEN "1110111111111111",
               x"D" WHEN "1101111111111111",
               x"E" WHEN "1011111111111111",
               x"F" WHEN "0111111111111111",
               x"0" WHEN OTHERS            ;


SliceDataOut   <= RdDataArray(Slv2Int(DecodedMiss));

END MainArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.CacheOutputDecoder(MainArch)
--PORT MAP   (Miss         => SLV,
--            RdDataArray  => SLV,
--            SliceDataOut => SLV
--           );
------------------------------------------------------------------------------------------