------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Project:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BasicPackage.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY MainMemoryTestbench IS
    
    PORT   (DataRd     : IN  uint32;
            Address    : IN  uint32;
            RdWrEnable : IN  uint02;
            DataWr     : OUT uint32 
           );
    
END ENTITY MainMemoryTestbench;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE TbArch OF MainMemoryTestbench IS

SIGNAL Tmp : uint32;

BEGIN

------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------

WITH RdWrEnable SELECT
DataWr <= Tmp         WHEN "10",
          Tmp         WHEN "11",
          x"FFFFFFFF" WHEN OTHERS;

WITH Address SELECT
Tmp    <= "00001111111111111111101010110111" WHEN (Int2Slv(000,32)),
          "00001111111111111111101010110111" WHEN (Int2Slv(000,32)),
          "01000000000000000000110110010011" WHEN (Int2Slv(001,32)),
          "00001011000000000000000001100111" WHEN (Int2Slv(002,32)),
          "00000001000000000000000001100111" WHEN (Int2Slv(016,32)),
          "00000010000000000000000001100111" WHEN (Int2Slv(032,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(033,32)),
          "00000000000010101010101000000011" WHEN (Int2Slv(048,32)),
          "00000000000100000000111110010011" WHEN (Int2Slv(049,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(050,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(051,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(052,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(053,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(054,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(055,32)),
          "00000000000000000000101000010011" WHEN (Int2Slv(064,32)),
          "00110000010011011010000001110011" WHEN (Int2Slv(065,32)),
          "00000000000000000000111110010011" WHEN (Int2Slv(066,32)),
          "00000000000100000000111100010011" WHEN (Int2Slv(067,32)),
          "00000000011000000000111010010011" WHEN (Int2Slv(068,32)),
          "00000000001000000000000010010011" WHEN (Int2Slv(069,32)),
          "00000000001100000000000100010011" WHEN (Int2Slv(070,32)),
          "00000000010000000000000110010011" WHEN (Int2Slv(071,32)),
          "00000000010100000000001000010011" WHEN (Int2Slv(072,32)),
          "00000000011000000000001010010011" WHEN (Int2Slv(073,32)),
          "00000000011100000000001100010011" WHEN (Int2Slv(074,32)),
          "00000000000100000000001110010011" WHEN (Int2Slv(075,32)),
          "00000000000000000000010110010011" WHEN (Int2Slv(076,32)),
          "00000000000000000000011000010011" WHEN (Int2Slv(077,32)),
          "00000000000000000000011010010011" WHEN (Int2Slv(078,32)),
          "00000000000000000000011100010011" WHEN (Int2Slv(079,32)),
          "00000000000000000000011110010011" WHEN (Int2Slv(080,32)),
          "00000000000000000000100000010011" WHEN (Int2Slv(081,32)),
          "00000000000110101000100010010011" WHEN (Int2Slv(082,32)),
          "00000001111011111000011101100011" WHEN (Int2Slv(083,32)),
          "00000101001000000000000001100111" WHEN (Int2Slv(084,32)),
          "00110000010011011011000001110011" WHEN (Int2Slv(096,32)),
          "00000000000110100101111000110011" WHEN (Int2Slv(097,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(098,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(099,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(100,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(101,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(102,32)),
          "00000001110111100000111000110011" WHEN (Int2Slv(103,32)),
          "00000010011100001000010110110011" WHEN (Int2Slv(104,32)),
          "00000010011100010000011000110011" WHEN (Int2Slv(105,32)),
          "00000010011100011000011010110011" WHEN (Int2Slv(106,32)),
          "00000010011100100000011100110011" WHEN (Int2Slv(107,32)),
          "00000010011100101000011110110011" WHEN (Int2Slv(108,32)),
          "00000010011100110000100000110011" WHEN (Int2Slv(109,32)),
          "00000000000100111000001110010011" WHEN (Int2Slv(110,32)),
          "00000001010001011001000111100011" WHEN (Int2Slv(111,32)),
          "00000000000110001010000000100011" WHEN (Int2Slv(112,32)),
          "00000000000110001000100010010011" WHEN (Int2Slv(113,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(114,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(115,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(116,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(117,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(118,32)),
          "00000001010001100001000111100011" WHEN (Int2Slv(119,32)),
          "00000000001010001010000000100011" WHEN (Int2Slv(120,32)),
          "00000000000110001000100010010011" WHEN (Int2Slv(121,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(122,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(123,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(124,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(125,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(126,32)),
          "00000001010001101001000111100011" WHEN (Int2Slv(127,32)),
          "00000000001110001010000000100011" WHEN (Int2Slv(128,32)),
          "00000000000110001000100010010011" WHEN (Int2Slv(129,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(130,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(131,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(132,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(133,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(134,32)),
          "00000001010001110001000111100011" WHEN (Int2Slv(135,32)),
          "00000000010010001010000000100011" WHEN (Int2Slv(136,32)),
          "00000000000110001000100010010011" WHEN (Int2Slv(137,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(138,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(139,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(140,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(141,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(142,32)),
          "00000001010001111001000111100011" WHEN (Int2Slv(143,32)),
          "00000000010110001010000000100011" WHEN (Int2Slv(144,32)),
          "00000000000110001000100010010011" WHEN (Int2Slv(145,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(146,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(147,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(148,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(149,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(150,32)),
          "00000001010010000001000111100011" WHEN (Int2Slv(151,32)),
          "00000000011010001010000000100011" WHEN (Int2Slv(152,32)),
          "00000000000110001000100010010011" WHEN (Int2Slv(153,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(154,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(155,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(156,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(157,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(158,32)),
          "11111110011111100101001111100011" WHEN (Int2Slv(159,32)),
          "00000000001000000000001110010011" WHEN (Int2Slv(160,32)),
          "00000001110100001000000010110011" WHEN (Int2Slv(161,32)),
          "00000001110100010000000100110011" WHEN (Int2Slv(162,32)),
          "00000001110100011000000110110011" WHEN (Int2Slv(163,32)),
          "00000001110100100000001000110011" WHEN (Int2Slv(164,32)),
          "00000001110100101000001010110011" WHEN (Int2Slv(165,32)),
          "00000001110100110000001100110011" WHEN (Int2Slv(166,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(167,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(168,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(169,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(170,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(171,32)),
          "11111100011011100101110101100011" WHEN (Int2Slv(172,32)),
          "00000101001000000000000001100111" WHEN (Int2Slv(173,32)),
          "11111111111111111111111111111111" WHEN OTHERS;
END TbArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.MainMemoryTestbench(TbArch)
--PORT MAP   (DataRd     => SLV,
--            Address    => SLV,
--            RdWrEnable => SLV,
--            DataWr     => SLV
--           );
------------------------------------------------------------------------------------------
