------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

USE WORK.BasicPackage.ALL;

ENTITY S2RegisterReadStageTestProtocol IS
END S2RegisterReadStageTestProtocol;

ARCHITECTURE S2RegisterReadStageTestProtocolArch OF S2RegisterReadStageTestProtocol IS

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------



BEGIN



END S2RegisterReadStageTestProtocolArch;
