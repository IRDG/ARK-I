------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

USE WORK.BasicPackage.ALL;

ENTITY S6ControlFsmTestProtocol IS
END S6ControlFsmTestProtocol;

ARCHITECTURE S6ControlFsmTestProtocolArch OF S6ControlFsmTestProtocol IS

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------



BEGIN



END S6ControlFsmTestProtocolArch;
