------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Proyect:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BasicPackage.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY Shifter IS
    
    PORT   (Input    : IN  uint32;
            Shamt    : IN  uint05;
            ArithRlN : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
            Output   : OUT uint32
           );
    
END ENTITY Shifter;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE MainArch OF Shifter IS

CONSTANT Zero           : STD_LOGIC := '0';

SIGNAL   ShiftLeftLogic : uint32;
SIGNAL   ShiftRghtLogic : uint32;
SIGNAL   ShiftRghtArith : uint32;

BEGIN

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

WITH ArithRlN SELECT
Output <= ShiftRghtLogic WHEN "00"  ,
          ShiftRghtArith WHEN "01"  ,
          ShiftLeftLogic WHEN "10"  ,
          ShiftLeftLogic WHEN OTHERS;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

WITH Shamt SELECT
ShiftLeftLogic( 0) <= Input( 0) WHEN "00000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 1) <= Input( 1) WHEN "00000",
                      Input( 0) WHEN "00001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 2) <= Input( 2) WHEN "00000",
                      Input( 1) WHEN "00001",
                      Input( 0) WHEN "00010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 3) <= Input( 3) WHEN "00000",
                      Input( 2) WHEN "00001",
                      Input( 1) WHEN "00010",
                      Input( 0) WHEN "00011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 4) <= Input( 4) WHEN "00000",
                      Input( 3) WHEN "00001",
                      Input( 2) WHEN "00010",
                      Input( 1) WHEN "00011",
                      Input( 0) WHEN "00100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 5) <= Input( 5) WHEN "00000",
                      Input( 4) WHEN "00001",
                      Input( 3) WHEN "00010",
                      Input( 2) WHEN "00011",
                      Input( 1) WHEN "00100",
                      Input( 0) WHEN "00101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 6) <= Input( 6) WHEN "00000",
                      Input( 5) WHEN "00001",
                      Input( 4) WHEN "00010",
                      Input( 3) WHEN "00011",
                      Input( 2) WHEN "00100",
                      Input( 1) WHEN "00101",
                      Input( 0) WHEN "00110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 7) <= Input( 7) WHEN "00000",
                      Input( 6) WHEN "00001",
                      Input( 5) WHEN "00010",
                      Input( 4) WHEN "00011",
                      Input( 3) WHEN "00100",
                      Input( 2) WHEN "00101",
                      Input( 1) WHEN "00110",
                      Input( 0) WHEN "00111",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 8) <= Input( 8) WHEN "00000",
                      Input( 7) WHEN "00001",
                      Input( 6) WHEN "00010",
                      Input( 5) WHEN "00011",
                      Input( 4) WHEN "00100",
                      Input( 3) WHEN "00101",
                      Input( 2) WHEN "00110",
                      Input( 1) WHEN "00111",
                      Input( 0) WHEN "01000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic( 9) <= Input( 9) WHEN "00000",
                      Input( 8) WHEN "00001",
                      Input( 7) WHEN "00010",
                      Input( 6) WHEN "00011",
                      Input( 5) WHEN "00100",
                      Input( 4) WHEN "00101",
                      Input( 3) WHEN "00110",
                      Input( 2) WHEN "00111",
                      Input( 1) WHEN "01000",
                      Input( 0) WHEN "01001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(10) <= Input(10) WHEN "00000",
                      Input( 9) WHEN "00001",
                      Input( 8) WHEN "00010",
                      Input( 7) WHEN "00011",
                      Input( 6) WHEN "00100",
                      Input( 5) WHEN "00101",
                      Input( 4) WHEN "00110",
                      Input( 3) WHEN "00111",
                      Input( 2) WHEN "01000",
                      Input( 1) WHEN "01001",
                      Input( 0) WHEN "01010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(11) <= Input(11) WHEN "00000",
                      Input(10) WHEN "00001",
                      Input( 9) WHEN "00010",
                      Input( 8) WHEN "00011",
                      Input( 7) WHEN "00100",
                      Input( 6) WHEN "00101",
                      Input( 5) WHEN "00110",
                      Input( 4) WHEN "00111",
                      Input( 3) WHEN "01000",
                      Input( 2) WHEN "01001",
                      Input( 1) WHEN "01010",
                      Input( 0) WHEN "01011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(12) <= Input(12) WHEN "00000",
                      Input(11) WHEN "00001",
                      Input(10) WHEN "00010",
                      Input( 9) WHEN "00011",
                      Input( 8) WHEN "00100",
                      Input( 7) WHEN "00101",
                      Input( 6) WHEN "00110",
                      Input( 5) WHEN "00111",
                      Input( 4) WHEN "01000",
                      Input( 3) WHEN "01001",
                      Input( 2) WHEN "01010",
                      Input( 1) WHEN "01011",
                      Input( 0) WHEN "01100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(13) <= Input(13) WHEN "00000",
                      Input(12) WHEN "00001",
                      Input(11) WHEN "00010",
                      Input(10) WHEN "00011",
                      Input( 9) WHEN "00100",
                      Input( 8) WHEN "00101",
                      Input( 7) WHEN "00110",
                      Input( 6) WHEN "00111",
                      Input( 5) WHEN "01000",
                      Input( 4) WHEN "01001",
                      Input( 3) WHEN "01010",
                      Input( 2) WHEN "01011",
                      Input( 1) WHEN "01100",
                      Input( 0) WHEN "01101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(14) <= Input(14) WHEN "00000",
                      Input(13) WHEN "00001",
                      Input(12) WHEN "00010",
                      Input(11) WHEN "00011",
                      Input(10) WHEN "00100",
                      Input( 9) WHEN "00101",
                      Input( 8) WHEN "00110",
                      Input( 7) WHEN "00111",
                      Input( 6) WHEN "01000",
                      Input( 5) WHEN "01001",
                      Input( 4) WHEN "01010",
                      Input( 3) WHEN "01011",
                      Input( 2) WHEN "01100",
                      Input( 1) WHEN "01101",
                      Input( 0) WHEN "01110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(15) <= Input(15) WHEN "00000",
                      Input(14) WHEN "00001",
                      Input(13) WHEN "00010",
                      Input(12) WHEN "00011",
                      Input(11) WHEN "00100",
                      Input(10) WHEN "00101",
                      Input( 9) WHEN "00110",
                      Input( 8) WHEN "00111",
                      Input( 7) WHEN "01000",
                      Input( 6) WHEN "01001",
                      Input( 5) WHEN "01010",
                      Input( 4) WHEN "01011",
                      Input( 3) WHEN "01100",
                      Input( 2) WHEN "01101",
                      Input( 1) WHEN "01110",
                      Input( 0) WHEN "01111",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(16) <= Input(16) WHEN "00000",
                      Input(15) WHEN "00001",
                      Input(14) WHEN "00010",
                      Input(13) WHEN "00011",
                      Input(12) WHEN "00100",
                      Input(11) WHEN "00101",
                      Input(10) WHEN "00110",
                      Input( 9) WHEN "00111",
                      Input( 8) WHEN "01000",
                      Input( 7) WHEN "01001",
                      Input( 6) WHEN "01010",
                      Input( 5) WHEN "01011",
                      Input( 4) WHEN "01100",
                      Input( 3) WHEN "01101",
                      Input( 2) WHEN "01110",
                      Input( 1) WHEN "01111",
                      Input( 0) WHEN "10000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(17) <= Input(17) WHEN "00000",
                      Input(16) WHEN "00001",
                      Input(15) WHEN "00010",
                      Input(14) WHEN "00011",
                      Input(13) WHEN "00100",
                      Input(12) WHEN "00101",
                      Input(11) WHEN "00110",
                      Input(10) WHEN "00111",
                      Input( 9) WHEN "01000",
                      Input( 8) WHEN "01001",
                      Input( 7) WHEN "01010",
                      Input( 6) WHEN "01011",
                      Input( 5) WHEN "01100",
                      Input( 4) WHEN "01101",
                      Input( 3) WHEN "01110",
                      Input( 2) WHEN "01111",
                      Input( 1) WHEN "10000",
                      Input( 0) WHEN "10001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(18) <= Input(18) WHEN "00000",
                      Input(17) WHEN "00001",
                      Input(16) WHEN "00010",
                      Input(15) WHEN "00011",
                      Input(14) WHEN "00100",
                      Input(13) WHEN "00101",
                      Input(12) WHEN "00110",
                      Input(11) WHEN "00111",
                      Input(10) WHEN "01000",
                      Input( 9) WHEN "01001",
                      Input( 8) WHEN "01010",
                      Input( 7) WHEN "01011",
                      Input( 6) WHEN "01100",
                      Input( 5) WHEN "01101",
                      Input( 4) WHEN "01110",
                      Input( 3) WHEN "01111",
                      Input( 2) WHEN "10000",
                      Input( 1) WHEN "10001",
                      Input( 0) WHEN "10010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(19) <= Input(19) WHEN "00000",
                      Input(18) WHEN "00001",
                      Input(17) WHEN "00010",
                      Input(16) WHEN "00011",
                      Input(15) WHEN "00100",
                      Input(14) WHEN "00101",
                      Input(13) WHEN "00110",
                      Input(12) WHEN "00111",
                      Input(11) WHEN "01000",
                      Input(10) WHEN "01001",
                      Input( 9) WHEN "01010",
                      Input( 8) WHEN "01011",
                      Input( 7) WHEN "01100",
                      Input( 6) WHEN "01101",
                      Input( 5) WHEN "01110",
                      Input( 4) WHEN "01111",
                      Input( 3) WHEN "10000",
                      Input( 2) WHEN "10001",
                      Input( 1) WHEN "10010",
                      Input( 0) WHEN "10011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(20) <= Input(20) WHEN "00000",
                      Input(19) WHEN "00001",
                      Input(18) WHEN "00010",
                      Input(17) WHEN "00011",
                      Input(16) WHEN "00100",
                      Input(15) WHEN "00101",
                      Input(14) WHEN "00110",
                      Input(13) WHEN "00111",
                      Input(12) WHEN "01000",
                      Input(11) WHEN "01001",
                      Input(10) WHEN "01010",
                      Input( 9) WHEN "01011",
                      Input( 8) WHEN "01100",
                      Input( 7) WHEN "01101",
                      Input( 6) WHEN "01110",
                      Input( 5) WHEN "01111",
                      Input( 4) WHEN "10000",
                      Input( 3) WHEN "10001",
                      Input( 2) WHEN "10010",
                      Input( 1) WHEN "10011",
                      Input( 0) WHEN "10100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(21) <= Input(21) WHEN "00000",
                      Input(20) WHEN "00001",
                      Input(19) WHEN "00010",
                      Input(18) WHEN "00011",
                      Input(17) WHEN "00100",
                      Input(16) WHEN "00101",
                      Input(15) WHEN "00110",
                      Input(14) WHEN "00111",
                      Input(13) WHEN "01000",
                      Input(12) WHEN "01001",
                      Input(11) WHEN "01010",
                      Input(10) WHEN "01011",
                      Input( 9) WHEN "01100",
                      Input( 8) WHEN "01101",
                      Input( 7) WHEN "01110",
                      Input( 6) WHEN "01111",
                      Input( 5) WHEN "10000",
                      Input( 4) WHEN "10001",
                      Input( 3) WHEN "10010",
                      Input( 2) WHEN "10011",
                      Input( 1) WHEN "10100",
                      Input( 0) WHEN "10101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(22) <= Input(22) WHEN "00000",
                      Input(21) WHEN "00001",
                      Input(20) WHEN "00010",
                      Input(19) WHEN "00011",
                      Input(18) WHEN "00100",
                      Input(17) WHEN "00101",
                      Input(16) WHEN "00110",
                      Input(15) WHEN "00111",
                      Input(14) WHEN "01000",
                      Input(13) WHEN "01001",
                      Input(12) WHEN "01010",
                      Input(11) WHEN "01011",
                      Input(10) WHEN "01100",
                      Input( 9) WHEN "01101",
                      Input( 8) WHEN "01110",
                      Input( 7) WHEN "01111",
                      Input( 6) WHEN "10000",
                      Input( 5) WHEN "10001",
                      Input( 4) WHEN "10010",
                      Input( 3) WHEN "10011",
                      Input( 2) WHEN "10100",
                      Input( 1) WHEN "10101",
                      Input( 0) WHEN "10110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(23) <= Input(23) WHEN "00000",
                      Input(22) WHEN "00001",
                      Input(21) WHEN "00010",
                      Input(20) WHEN "00011",
                      Input(19) WHEN "00100",
                      Input(18) WHEN "00101",
                      Input(17) WHEN "00110",
                      Input(16) WHEN "00111",
                      Input(15) WHEN "01000",
                      Input(14) WHEN "01001",
                      Input(13) WHEN "01010",
                      Input(12) WHEN "01011",
                      Input(11) WHEN "01100",
                      Input(10) WHEN "01101",
                      Input( 9) WHEN "01110",
                      Input( 8) WHEN "01111",
                      Input( 7) WHEN "10000",
                      Input( 6) WHEN "10001",
                      Input( 5) WHEN "10010",
                      Input( 4) WHEN "10011",
                      Input( 3) WHEN "10100",
                      Input( 2) WHEN "10101",
                      Input( 1) WHEN "10110",
                      Input( 0) WHEN "10111",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(24) <= Input(24) WHEN "00000",
                      Input(23) WHEN "00001",
                      Input(22) WHEN "00010",
                      Input(21) WHEN "00011",
                      Input(20) WHEN "00100",
                      Input(19) WHEN "00101",
                      Input(18) WHEN "00110",
                      Input(17) WHEN "00111",
                      Input(16) WHEN "01000",
                      Input(15) WHEN "01001",
                      Input(14) WHEN "01010",
                      Input(13) WHEN "01011",
                      Input(12) WHEN "01100",
                      Input(11) WHEN "01101",
                      Input(10) WHEN "01110",
                      Input( 9) WHEN "01111",
                      Input( 8) WHEN "10000",
                      Input( 7) WHEN "10001",
                      Input( 6) WHEN "10010",
                      Input( 5) WHEN "10011",
                      Input( 4) WHEN "10100",
                      Input( 3) WHEN "10101",
                      Input( 2) WHEN "10110",
                      Input( 1) WHEN "10111",
                      Input( 0) WHEN "11000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(25) <= Input(25) WHEN "00000",
                      Input(24) WHEN "00001",
                      Input(23) WHEN "00010",
                      Input(22) WHEN "00011",
                      Input(21) WHEN "00100",
                      Input(20) WHEN "00101",
                      Input(19) WHEN "00110",
                      Input(18) WHEN "00111",
                      Input(17) WHEN "01000",
                      Input(16) WHEN "01001",
                      Input(15) WHEN "01010",
                      Input(14) WHEN "01011",
                      Input(13) WHEN "01100",
                      Input(12) WHEN "01101",
                      Input(11) WHEN "01110",
                      Input(10) WHEN "01111",
                      Input( 9) WHEN "10000",
                      Input( 8) WHEN "10001",
                      Input( 7) WHEN "10010",
                      Input( 6) WHEN "10011",
                      Input( 5) WHEN "10100",
                      Input( 4) WHEN "10101",
                      Input( 3) WHEN "10110",
                      Input( 2) WHEN "10111",
                      Input( 1) WHEN "11000",
                      Input( 0) WHEN "11001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(26) <= Input(26) WHEN "00000",
                      Input(25) WHEN "00001",
                      Input(24) WHEN "00010",
                      Input(23) WHEN "00011",
                      Input(22) WHEN "00100",
                      Input(21) WHEN "00101",
                      Input(20) WHEN "00110",
                      Input(19) WHEN "00111",
                      Input(18) WHEN "01000",
                      Input(17) WHEN "01001",
                      Input(16) WHEN "01010",
                      Input(15) WHEN "01011",
                      Input(14) WHEN "01100",
                      Input(13) WHEN "01101",
                      Input(12) WHEN "01110",
                      Input(11) WHEN "01111",
                      Input(10) WHEN "10000",
                      Input( 9) WHEN "10001",
                      Input( 8) WHEN "10010",
                      Input( 7) WHEN "10011",
                      Input( 6) WHEN "10100",
                      Input( 5) WHEN "10101",
                      Input( 4) WHEN "10110",
                      Input( 3) WHEN "10111",
                      Input( 2) WHEN "11000",
                      Input( 1) WHEN "11001",
                      Input( 0) WHEN "11010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(27) <= Input(27) WHEN "00000",
                      Input(26) WHEN "00001",
                      Input(25) WHEN "00010",
                      Input(24) WHEN "00011",
                      Input(23) WHEN "00100",
                      Input(22) WHEN "00101",
                      Input(21) WHEN "00110",
                      Input(20) WHEN "00111",
                      Input(19) WHEN "01000",
                      Input(18) WHEN "01001",
                      Input(17) WHEN "01010",
                      Input(16) WHEN "01011",
                      Input(15) WHEN "01100",
                      Input(14) WHEN "01101",
                      Input(13) WHEN "01110",
                      Input(12) WHEN "01111",
                      Input(11) WHEN "10000",
                      Input(10) WHEN "10001",
                      Input( 9) WHEN "10010",
                      Input( 8) WHEN "10011",
                      Input( 7) WHEN "10100",
                      Input( 6) WHEN "10101",
                      Input( 5) WHEN "10110",
                      Input( 4) WHEN "10111",
                      Input( 3) WHEN "11000",
                      Input( 2) WHEN "11001",
                      Input( 1) WHEN "11010",
                      Input( 0) WHEN "11011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(28) <= Input(28) WHEN "00000",
                      Input(27) WHEN "00001",
                      Input(26) WHEN "00010",
                      Input(25) WHEN "00011",
                      Input(24) WHEN "00100",
                      Input(23) WHEN "00101",
                      Input(22) WHEN "00110",
                      Input(21) WHEN "00111",
                      Input(20) WHEN "01000",
                      Input(19) WHEN "01001",
                      Input(18) WHEN "01010",
                      Input(17) WHEN "01011",
                      Input(16) WHEN "01100",
                      Input(15) WHEN "01101",
                      Input(14) WHEN "01110",
                      Input(13) WHEN "01111",
                      Input(12) WHEN "10000",
                      Input(11) WHEN "10001",
                      Input(10) WHEN "10010",
                      Input( 9) WHEN "10011",
                      Input( 8) WHEN "10100",
                      Input( 7) WHEN "10101",
                      Input( 6) WHEN "10110",
                      Input( 5) WHEN "10111",
                      Input( 4) WHEN "11000",
                      Input( 3) WHEN "11001",
                      Input( 2) WHEN "11010",
                      Input( 1) WHEN "11011",
                      Input( 0) WHEN "11100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(29) <= Input(29) WHEN "00000",
                      Input(28) WHEN "00001",
                      Input(27) WHEN "00010",
                      Input(26) WHEN "00011",
                      Input(25) WHEN "00100",
                      Input(24) WHEN "00101",
                      Input(23) WHEN "00110",
                      Input(22) WHEN "00111",
                      Input(21) WHEN "01000",
                      Input(20) WHEN "01001",
                      Input(19) WHEN "01010",
                      Input(18) WHEN "01011",
                      Input(17) WHEN "01100",
                      Input(16) WHEN "01101",
                      Input(15) WHEN "01110",
                      Input(14) WHEN "01111",
                      Input(13) WHEN "10000",
                      Input(12) WHEN "10001",
                      Input(11) WHEN "10010",
                      Input(10) WHEN "10011",
                      Input( 9) WHEN "10100",
                      Input( 8) WHEN "10101",
                      Input( 7) WHEN "10110",
                      Input( 6) WHEN "10111",
                      Input( 5) WHEN "11000",
                      Input( 4) WHEN "11001",
                      Input( 3) WHEN "11010",
                      Input( 2) WHEN "11011",
                      Input( 1) WHEN "11100",
                      Input( 0) WHEN "11101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(30) <= Input(30) WHEN "00000",
                      Input(29) WHEN "00001",
                      Input(28) WHEN "00010",
                      Input(27) WHEN "00011",
                      Input(26) WHEN "00100",
                      Input(25) WHEN "00101",
                      Input(24) WHEN "00110",
                      Input(23) WHEN "00111",
                      Input(22) WHEN "01000",
                      Input(21) WHEN "01001",
                      Input(20) WHEN "01010",
                      Input(19) WHEN "01011",
                      Input(18) WHEN "01100",
                      Input(17) WHEN "01101",
                      Input(16) WHEN "01110",
                      Input(15) WHEN "01111",
                      Input(14) WHEN "10000",
                      Input(13) WHEN "10001",
                      Input(12) WHEN "10010",
                      Input(11) WHEN "10011",
                      Input(10) WHEN "10100",
                      Input( 9) WHEN "10101",
                      Input( 8) WHEN "10110",
                      Input( 7) WHEN "10111",
                      Input( 6) WHEN "11000",
                      Input( 5) WHEN "11001",
                      Input( 4) WHEN "11010",
                      Input( 3) WHEN "11011",
                      Input( 2) WHEN "11100",
                      Input( 1) WHEN "11101",
                      Input( 0) WHEN "11110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftLeftLogic(31) <= Input(31) WHEN "00000",
                      Input(30) WHEN "00001",
                      Input(29) WHEN "00010",
                      Input(28) WHEN "00011",
                      Input(27) WHEN "00100",
                      Input(26) WHEN "00101",
                      Input(25) WHEN "00110",
                      Input(24) WHEN "00111",
                      Input(23) WHEN "01000",
                      Input(22) WHEN "01001",
                      Input(21) WHEN "01010",
                      Input(20) WHEN "01011",
                      Input(19) WHEN "01100",
                      Input(18) WHEN "01101",
                      Input(17) WHEN "01110",
                      Input(16) WHEN "01111",
                      Input(15) WHEN "10000",
                      Input(14) WHEN "10001",
                      Input(13) WHEN "10010",
                      Input(12) WHEN "10011",
                      Input(11) WHEN "10100",
                      Input(10) WHEN "10101",
                      Input( 9) WHEN "10110",
                      Input( 8) WHEN "10111",
                      Input( 7) WHEN "11000",
                      Input( 6) WHEN "11001",
                      Input( 5) WHEN "11010",
                      Input( 4) WHEN "11011",
                      Input( 3) WHEN "11100",
                      Input( 2) WHEN "11101",
                      Input( 1) WHEN "11110",
                      Input( 0) WHEN "11111",
                      Zero      WHEN OTHERS ;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

WITH Shamt SELECT
ShiftRghtLogic( 0) <= Input( 0) WHEN "00000",
                      Input( 1) WHEN "00001",
                      Input( 2) WHEN "00010",
                      Input( 3) WHEN "00011",
                      Input( 4) WHEN "00100",
                      Input( 5) WHEN "00101",
                      Input( 6) WHEN "00110",
                      Input( 7) WHEN "00111",
                      Input( 8) WHEN "01000",
                      Input( 9) WHEN "01001",
                      Input(10) WHEN "01010",
                      Input(11) WHEN "01011",
                      Input(12) WHEN "01100",
                      Input(13) WHEN "01101",
                      Input(14) WHEN "01110",
                      Input(15) WHEN "01111",
                      Input(16) WHEN "10000",
                      Input(17) WHEN "10001",
                      Input(18) WHEN "10010",
                      Input(19) WHEN "10011",
                      Input(20) WHEN "10100",
                      Input(21) WHEN "10101",
                      Input(22) WHEN "10110",
                      Input(23) WHEN "10111",
                      Input(24) WHEN "11000",
                      Input(25) WHEN "11001",
                      Input(26) WHEN "11010",
                      Input(27) WHEN "11011",
                      Input(28) WHEN "11100",
                      Input(29) WHEN "11101",
                      Input(30) WHEN "11110",
                      Input(31) WHEN OTHERS ;
                      
WITH Shamt SELECT
ShiftRghtLogic( 1) <= Input( 1) WHEN "00000",
                      Input( 2) WHEN "00001",
                      Input( 3) WHEN "00010",
                      Input( 4) WHEN "00011",
                      Input( 5) WHEN "00100",
                      Input( 6) WHEN "00101",
                      Input( 7) WHEN "00110",
                      Input( 8) WHEN "00111",
                      Input( 9) WHEN "01000",
                      Input(10) WHEN "01001",
                      Input(11) WHEN "01010",
                      Input(12) WHEN "01011",
                      Input(13) WHEN "01100",
                      Input(14) WHEN "01101",
                      Input(15) WHEN "01110",
                      Input(16) WHEN "01111",
                      Input(17) WHEN "10000",
                      Input(18) WHEN "10001",
                      Input(19) WHEN "10010",
                      Input(20) WHEN "10011",
                      Input(21) WHEN "10100",
                      Input(22) WHEN "10101",
                      Input(23) WHEN "10110",
                      Input(24) WHEN "10111",
                      Input(25) WHEN "11000",
                      Input(26) WHEN "11001",
                      Input(27) WHEN "11010",
                      Input(28) WHEN "11011",
                      Input(29) WHEN "11100",
                      Input(30) WHEN "11101",
                      Input(31) WHEN "11110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 2) <= Input( 2) WHEN "00000",
                      Input( 3) WHEN "00001",
                      Input( 4) WHEN "00010",
                      Input( 5) WHEN "00011",
                      Input( 6) WHEN "00100",
                      Input( 7) WHEN "00101",
                      Input( 8) WHEN "00110",
                      Input( 9) WHEN "00111",
                      Input(10) WHEN "01000",
                      Input(11) WHEN "01001",
                      Input(12) WHEN "01010",
                      Input(13) WHEN "01011",
                      Input(14) WHEN "01100",
                      Input(15) WHEN "01101",
                      Input(16) WHEN "01110",
                      Input(17) WHEN "01111",
                      Input(18) WHEN "10000",
                      Input(19) WHEN "10001",
                      Input(20) WHEN "10010",
                      Input(21) WHEN "10011",
                      Input(22) WHEN "10100",
                      Input(23) WHEN "10101",
                      Input(24) WHEN "10110",
                      Input(25) WHEN "10111",
                      Input(26) WHEN "11000",
                      Input(27) WHEN "11001",
                      Input(28) WHEN "11010",
                      Input(29) WHEN "11011",
                      Input(30) WHEN "11100",
                      Input(31) WHEN "11101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 3) <= Input( 3) WHEN "00000",
                      Input( 4) WHEN "00001",
                      Input( 5) WHEN "00010",
                      Input( 6) WHEN "00011",
                      Input( 7) WHEN "00100",
                      Input( 8) WHEN "00101",
                      Input( 9) WHEN "00110",
                      Input(10) WHEN "00111",
                      Input(11) WHEN "01000",
                      Input(12) WHEN "01001",
                      Input(13) WHEN "01010",
                      Input(14) WHEN "01011",
                      Input(15) WHEN "01100",
                      Input(16) WHEN "01101",
                      Input(17) WHEN "01110",
                      Input(18) WHEN "01111",
                      Input(19) WHEN "10000",
                      Input(20) WHEN "10001",
                      Input(21) WHEN "10010",
                      Input(22) WHEN "10011",
                      Input(23) WHEN "10100",
                      Input(24) WHEN "10101",
                      Input(25) WHEN "10110",
                      Input(26) WHEN "10111",
                      Input(27) WHEN "11000",
                      Input(28) WHEN "11001",
                      Input(29) WHEN "11010",
                      Input(30) WHEN "11011",
                      Input(31) WHEN "11100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 4) <= Input( 4) WHEN "00000",
                      Input( 5) WHEN "00001",
                      Input( 6) WHEN "00010",
                      Input( 7) WHEN "00011",
                      Input( 8) WHEN "00100",
                      Input( 9) WHEN "00101",
                      Input(10) WHEN "00110",
                      Input(11) WHEN "00111",
                      Input(12) WHEN "01000",
                      Input(13) WHEN "01001",
                      Input(14) WHEN "01010",
                      Input(15) WHEN "01011",
                      Input(16) WHEN "01100",
                      Input(17) WHEN "01101",
                      Input(18) WHEN "01110",
                      Input(19) WHEN "01111",
                      Input(20) WHEN "10000",
                      Input(21) WHEN "10001",
                      Input(22) WHEN "10010",
                      Input(23) WHEN "10011",
                      Input(24) WHEN "10100",
                      Input(25) WHEN "10101",
                      Input(26) WHEN "10110",
                      Input(27) WHEN "10111",
                      Input(28) WHEN "11000",
                      Input(29) WHEN "11001",
                      Input(30) WHEN "11010",
                      Input(31) WHEN "11011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 5) <= Input( 5) WHEN "00000",
                      Input( 6) WHEN "00001",
                      Input( 7) WHEN "00010",
                      Input( 8) WHEN "00011",
                      Input( 9) WHEN "00100",
                      Input(10) WHEN "00101",
                      Input(11) WHEN "00110",
                      Input(12) WHEN "00111",
                      Input(13) WHEN "01000",
                      Input(14) WHEN "01001",
                      Input(15) WHEN "01010",
                      Input(16) WHEN "01011",
                      Input(17) WHEN "01100",
                      Input(18) WHEN "01101",
                      Input(19) WHEN "01110",
                      Input(20) WHEN "01111",
                      Input(21) WHEN "10000",
                      Input(22) WHEN "10001",
                      Input(23) WHEN "10010",
                      Input(24) WHEN "10011",
                      Input(25) WHEN "10100",
                      Input(26) WHEN "10101",
                      Input(27) WHEN "10110",
                      Input(28) WHEN "10111",
                      Input(29) WHEN "11000",
                      Input(30) WHEN "11001",
                      Input(31) WHEN "11010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 6) <= Input( 6) WHEN "00000",
                      Input( 7) WHEN "00001",
                      Input( 8) WHEN "00010",
                      Input( 9) WHEN "00011",
                      Input(10) WHEN "00100",
                      Input(11) WHEN "00101",
                      Input(12) WHEN "00110",
                      Input(13) WHEN "00111",
                      Input(14) WHEN "01000",
                      Input(15) WHEN "01001",
                      Input(16) WHEN "01010",
                      Input(17) WHEN "01011",
                      Input(18) WHEN "01100",
                      Input(19) WHEN "01101",
                      Input(20) WHEN "01110",
                      Input(21) WHEN "01111",
                      Input(22) WHEN "10000",
                      Input(23) WHEN "10001",
                      Input(24) WHEN "10010",
                      Input(25) WHEN "10011",
                      Input(26) WHEN "10100",
                      Input(27) WHEN "10101",
                      Input(28) WHEN "10110",
                      Input(29) WHEN "10111",
                      Input(30) WHEN "11000",
                      Input(31) WHEN "11001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 7) <= Input( 7) WHEN "00000",
                      Input( 8) WHEN "00001",
                      Input( 9) WHEN "00010",
                      Input(10) WHEN "00011",
                      Input(11) WHEN "00100",
                      Input(12) WHEN "00101",
                      Input(13) WHEN "00110",
                      Input(14) WHEN "00111",
                      Input(15) WHEN "01000",
                      Input(16) WHEN "01001",
                      Input(17) WHEN "01010",
                      Input(18) WHEN "01011",
                      Input(19) WHEN "01100",
                      Input(20) WHEN "01101",
                      Input(21) WHEN "01110",
                      Input(22) WHEN "01111",
                      Input(23) WHEN "10000",
                      Input(24) WHEN "10001",
                      Input(25) WHEN "10010",
                      Input(26) WHEN "10011",
                      Input(27) WHEN "10100",
                      Input(28) WHEN "10101",
                      Input(29) WHEN "10110",
                      Input(30) WHEN "10111",
                      Input(31) WHEN "11000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 8) <= Input( 8) WHEN "00000",
                      Input( 9) WHEN "00001",
                      Input(10) WHEN "00010",
                      Input(11) WHEN "00011",
                      Input(12) WHEN "00100",
                      Input(13) WHEN "00101",
                      Input(14) WHEN "00110",
                      Input(15) WHEN "00111",
                      Input(16) WHEN "01000",
                      Input(17) WHEN "01001",
                      Input(18) WHEN "01010",
                      Input(19) WHEN "01011",
                      Input(20) WHEN "01100",
                      Input(21) WHEN "01101",
                      Input(22) WHEN "01110",
                      Input(23) WHEN "01111",
                      Input(24) WHEN "10000",
                      Input(25) WHEN "10001",
                      Input(26) WHEN "10010",
                      Input(27) WHEN "10011",
                      Input(28) WHEN "10100",
                      Input(29) WHEN "10101",
                      Input(30) WHEN "10110",
                      Input(31) WHEN "10111",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic( 9) <= Input( 9) WHEN "00000",
                      Input(10) WHEN "00001",
                      Input(11) WHEN "00010",
                      Input(12) WHEN "00011",
                      Input(13) WHEN "00100",
                      Input(14) WHEN "00101",
                      Input(15) WHEN "00110",
                      Input(16) WHEN "00111",
                      Input(17) WHEN "01000",
                      Input(18) WHEN "01001",
                      Input(19) WHEN "01010",
                      Input(20) WHEN "01011",
                      Input(21) WHEN "01100",
                      Input(22) WHEN "01101",
                      Input(23) WHEN "01110",
                      Input(24) WHEN "01111",
                      Input(25) WHEN "10000",
                      Input(26) WHEN "10001",
                      Input(27) WHEN "10010",
                      Input(28) WHEN "10011",
                      Input(29) WHEN "10100",
                      Input(30) WHEN "10101",
                      Input(31) WHEN "10110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(10) <= Input(10) WHEN "00000",
                      Input(11) WHEN "00001",
                      Input(12) WHEN "00010",
                      Input(13) WHEN "00011",
                      Input(14) WHEN "00100",
                      Input(15) WHEN "00101",
                      Input(16) WHEN "00110",
                      Input(17) WHEN "00111",
                      Input(18) WHEN "01000",
                      Input(19) WHEN "01001",
                      Input(20) WHEN "01010",
                      Input(21) WHEN "01011",
                      Input(22) WHEN "01100",
                      Input(23) WHEN "01101",
                      Input(24) WHEN "01110",
                      Input(25) WHEN "01111",
                      Input(26) WHEN "10000",
                      Input(27) WHEN "10001",
                      Input(28) WHEN "10010",
                      Input(29) WHEN "10011",
                      Input(30) WHEN "10100",
                      Input(31) WHEN "10101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(11) <= Input(11) WHEN "00000",
                      Input(12) WHEN "00001",
                      Input(13) WHEN "00010",
                      Input(14) WHEN "00011",
                      Input(15) WHEN "00100",
                      Input(16) WHEN "00101",
                      Input(17) WHEN "00110",
                      Input(18) WHEN "00111",
                      Input(19) WHEN "01000",
                      Input(20) WHEN "01001",
                      Input(21) WHEN "01010",
                      Input(22) WHEN "01011",
                      Input(23) WHEN "01100",
                      Input(24) WHEN "01101",
                      Input(25) WHEN "01110",
                      Input(26) WHEN "01111",
                      Input(27) WHEN "10000",
                      Input(28) WHEN "10001",
                      Input(29) WHEN "10010",
                      Input(30) WHEN "10011",
                      Input(31) WHEN "10100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(12) <= Input(12) WHEN "00000",
                      Input(13) WHEN "00001",
                      Input(14) WHEN "00010",
                      Input(15) WHEN "00011",
                      Input(16) WHEN "00100",
                      Input(17) WHEN "00101",
                      Input(18) WHEN "00110",
                      Input(19) WHEN "00111",
                      Input(20) WHEN "01000",
                      Input(21) WHEN "01001",
                      Input(22) WHEN "01010",
                      Input(23) WHEN "01011",
                      Input(24) WHEN "01100",
                      Input(25) WHEN "01101",
                      Input(26) WHEN "01110",
                      Input(27) WHEN "01111",
                      Input(28) WHEN "10000",
                      Input(29) WHEN "10001",
                      Input(30) WHEN "10010",
                      Input(31) WHEN "10011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(13) <= Input(13) WHEN "00000",
                      Input(14) WHEN "00001",
                      Input(15) WHEN "00010",
                      Input(16) WHEN "00011",
                      Input(17) WHEN "00100",
                      Input(18) WHEN "00101",
                      Input(19) WHEN "00110",
                      Input(20) WHEN "00111",
                      Input(21) WHEN "01000",
                      Input(22) WHEN "01001",
                      Input(23) WHEN "01010",
                      Input(24) WHEN "01011",
                      Input(25) WHEN "01100",
                      Input(26) WHEN "01101",
                      Input(27) WHEN "01110",
                      Input(28) WHEN "01111",
                      Input(29) WHEN "10000",
                      Input(30) WHEN "10001",
                      Input(31) WHEN "10010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(14) <= Input(14) WHEN "00000",
                      Input(15) WHEN "00001",
                      Input(16) WHEN "00010",
                      Input(17) WHEN "00011",
                      Input(18) WHEN "00100",
                      Input(19) WHEN "00101",
                      Input(20) WHEN "00110",
                      Input(21) WHEN "00111",
                      Input(22) WHEN "01000",
                      Input(23) WHEN "01001",
                      Input(24) WHEN "01010",
                      Input(25) WHEN "01011",
                      Input(26) WHEN "01100",
                      Input(27) WHEN "01101",
                      Input(28) WHEN "01110",
                      Input(29) WHEN "01111",
                      Input(30) WHEN "10000",
                      Input(31) WHEN "10001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(15) <= Input(15) WHEN "00000",
                      Input(16) WHEN "00001",
                      Input(17) WHEN "00010",
                      Input(18) WHEN "00011",
                      Input(19) WHEN "00100",
                      Input(20) WHEN "00101",
                      Input(21) WHEN "00110",
                      Input(22) WHEN "00111",
                      Input(23) WHEN "01000",
                      Input(24) WHEN "01001",
                      Input(25) WHEN "01010",
                      Input(26) WHEN "01011",
                      Input(27) WHEN "01100",
                      Input(28) WHEN "01101",
                      Input(29) WHEN "01110",
                      Input(30) WHEN "01111",
                      Input(31) WHEN "10000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(16) <= Input(16) WHEN "00000",
                      Input(17) WHEN "00001",
                      Input(18) WHEN "00010",
                      Input(19) WHEN "00011",
                      Input(20) WHEN "00100",
                      Input(21) WHEN "00101",
                      Input(22) WHEN "00110",
                      Input(23) WHEN "00111",
                      Input(24) WHEN "01000",
                      Input(25) WHEN "01001",
                      Input(26) WHEN "01010",
                      Input(27) WHEN "01011",
                      Input(28) WHEN "01100",
                      Input(29) WHEN "01101",
                      Input(30) WHEN "01110",
                      Input(31) WHEN "01111",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(17) <= Input(17) WHEN "00000",
                      Input(18) WHEN "00001",
                      Input(19) WHEN "00010",
                      Input(20) WHEN "00011",
                      Input(21) WHEN "00100",
                      Input(22) WHEN "00101",
                      Input(23) WHEN "00110",
                      Input(24) WHEN "00111",
                      Input(25) WHEN "01000",
                      Input(26) WHEN "01001",
                      Input(27) WHEN "01010",
                      Input(28) WHEN "01011",
                      Input(29) WHEN "01100",
                      Input(30) WHEN "01101",
                      Input(31) WHEN "01110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(18) <= Input(18) WHEN "00000",
                      Input(19) WHEN "00001",
                      Input(20) WHEN "00010",
                      Input(21) WHEN "00011",
                      Input(22) WHEN "00100",
                      Input(23) WHEN "00101",
                      Input(24) WHEN "00110",
                      Input(25) WHEN "00111",
                      Input(26) WHEN "01000",
                      Input(27) WHEN "01001",
                      Input(28) WHEN "01010",
                      Input(29) WHEN "01011",
                      Input(30) WHEN "01100",
                      Input(31) WHEN "01101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(19) <= Input(19) WHEN "00000",
                      Input(20) WHEN "00001",
                      Input(21) WHEN "00010",
                      Input(22) WHEN "00011",
                      Input(23) WHEN "00100",
                      Input(24) WHEN "00101",
                      Input(25) WHEN "00110",
                      Input(26) WHEN "00111",
                      Input(27) WHEN "01000",
                      Input(28) WHEN "01001",
                      Input(29) WHEN "01010",
                      Input(30) WHEN "01011",
                      Input(31) WHEN "01100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(20) <= Input(20) WHEN "00000",
                      Input(21) WHEN "00001",
                      Input(22) WHEN "00010",
                      Input(23) WHEN "00011",
                      Input(24) WHEN "00100",
                      Input(25) WHEN "00101",
                      Input(26) WHEN "00110",
                      Input(27) WHEN "00111",
                      Input(28) WHEN "01000",
                      Input(29) WHEN "01001",
                      Input(30) WHEN "01010",
                      Input(31) WHEN "01011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(21) <= Input(21) WHEN "00000",
                      Input(22) WHEN "00001",
                      Input(23) WHEN "00010",
                      Input(24) WHEN "00011",
                      Input(25) WHEN "00100",
                      Input(26) WHEN "00101",
                      Input(27) WHEN "00110",
                      Input(28) WHEN "00111",
                      Input(29) WHEN "01000",
                      Input(30) WHEN "01001",
                      Input(31) WHEN "01010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(22) <= Input(22) WHEN "00000",
                      Input(23) WHEN "00001",
                      Input(24) WHEN "00010",
                      Input(25) WHEN "00011",
                      Input(26) WHEN "00100",
                      Input(27) WHEN "00101",
                      Input(28) WHEN "00110",
                      Input(29) WHEN "00111",
                      Input(30) WHEN "01000",
                      Input(31) WHEN "01001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(23) <= Input(23) WHEN "00000",
                      Input(24) WHEN "00001",
                      Input(25) WHEN "00010",
                      Input(26) WHEN "00011",
                      Input(27) WHEN "00100",
                      Input(28) WHEN "00101",
                      Input(29) WHEN "00110",
                      Input(30) WHEN "00111",
                      Input(31) WHEN "01000",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(24) <= Input(24) WHEN "00000",
                      Input(25) WHEN "00001",
                      Input(26) WHEN "00010",
                      Input(27) WHEN "00011",
                      Input(28) WHEN "00100",
                      Input(29) WHEN "00101",
                      Input(30) WHEN "00110",
                      Input(31) WHEN "00111",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(25) <= Input(25) WHEN "00000",
                      Input(26) WHEN "00001",
                      Input(27) WHEN "00010",
                      Input(28) WHEN "00011",
                      Input(29) WHEN "00100",
                      Input(30) WHEN "00101",
                      Input(31) WHEN "00110",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(26) <= Input(26) WHEN "00000",
                      Input(27) WHEN "00001",
                      Input(28) WHEN "00010",
                      Input(29) WHEN "00011",
                      Input(30) WHEN "00100",
                      Input(31) WHEN "00101",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(27) <= Input(27) WHEN "00000",
                      Input(28) WHEN "00001",
                      Input(29) WHEN "00010",
                      Input(30) WHEN "00011",
                      Input(31) WHEN "00100",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(28) <= Input(28) WHEN "00000",
                      Input(29) WHEN "00001",
                      Input(30) WHEN "00010",
                      Input(31) WHEN "00011",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(29) <= Input(29) WHEN "00000",
                      Input(30) WHEN "00001",
                      Input(31) WHEN "00010",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(30) <= Input(30) WHEN "00000",
                      Input(31) WHEN "00001",
                      Zero      WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtLogic(31) <= Input(31) WHEN "00000",
                      Zero      WHEN OTHERS ;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

WITH Shamt SELECT
ShiftRghtArith( 0) <= Input( 0) WHEN "00000",
                      Input( 1) WHEN "00001",
                      Input( 2) WHEN "00010",
                      Input( 3) WHEN "00011",
                      Input( 4) WHEN "00100",
                      Input( 5) WHEN "00101",
                      Input( 6) WHEN "00110",
                      Input( 7) WHEN "00111",
                      Input( 8) WHEN "01000",
                      Input( 9) WHEN "01001",
                      Input(10) WHEN "01010",
                      Input(11) WHEN "01011",
                      Input(12) WHEN "01100",
                      Input(13) WHEN "01101",
                      Input(14) WHEN "01110",
                      Input(15) WHEN "01111",
                      Input(16) WHEN "10000",
                      Input(17) WHEN "10001",
                      Input(18) WHEN "10010",
                      Input(19) WHEN "10011",
                      Input(20) WHEN "10100",
                      Input(21) WHEN "10101",
                      Input(22) WHEN "10110",
                      Input(23) WHEN "10111",
                      Input(24) WHEN "11000",
                      Input(25) WHEN "11001",
                      Input(26) WHEN "11010",
                      Input(27) WHEN "11011",
                      Input(28) WHEN "11100",
                      Input(29) WHEN "11101",
                      Input(30) WHEN "11110",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 1) <= Input( 1) WHEN "00000",
                      Input( 2) WHEN "00001",
                      Input( 3) WHEN "00010",
                      Input( 4) WHEN "00011",
                      Input( 5) WHEN "00100",
                      Input( 6) WHEN "00101",
                      Input( 7) WHEN "00110",
                      Input( 8) WHEN "00111",
                      Input( 9) WHEN "01000",
                      Input(10) WHEN "01001",
                      Input(11) WHEN "01010",
                      Input(12) WHEN "01011",
                      Input(13) WHEN "01100",
                      Input(14) WHEN "01101",
                      Input(15) WHEN "01110",
                      Input(16) WHEN "01111",
                      Input(17) WHEN "10000",
                      Input(18) WHEN "10001",
                      Input(19) WHEN "10010",
                      Input(20) WHEN "10011",
                      Input(21) WHEN "10100",
                      Input(22) WHEN "10101",
                      Input(23) WHEN "10110",
                      Input(24) WHEN "10111",
                      Input(25) WHEN "11000",
                      Input(26) WHEN "11001",
                      Input(27) WHEN "11010",
                      Input(28) WHEN "11011",
                      Input(29) WHEN "11100",
                      Input(30) WHEN "11101",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 2) <= Input( 2) WHEN "00000",
                      Input( 3) WHEN "00001",
                      Input( 4) WHEN "00010",
                      Input( 5) WHEN "00011",
                      Input( 6) WHEN "00100",
                      Input( 7) WHEN "00101",
                      Input( 8) WHEN "00110",
                      Input( 9) WHEN "00111",
                      Input(10) WHEN "01000",
                      Input(11) WHEN "01001",
                      Input(12) WHEN "01010",
                      Input(13) WHEN "01011",
                      Input(14) WHEN "01100",
                      Input(15) WHEN "01101",
                      Input(16) WHEN "01110",
                      Input(17) WHEN "01111",
                      Input(18) WHEN "10000",
                      Input(19) WHEN "10001",
                      Input(20) WHEN "10010",
                      Input(21) WHEN "10011",
                      Input(22) WHEN "10100",
                      Input(23) WHEN "10101",
                      Input(24) WHEN "10110",
                      Input(25) WHEN "10111",
                      Input(26) WHEN "11000",
                      Input(27) WHEN "11001",
                      Input(28) WHEN "11010",
                      Input(29) WHEN "11011",
                      Input(30) WHEN "11100",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 3) <= Input( 3) WHEN "00000",
                      Input( 4) WHEN "00001",
                      Input( 5) WHEN "00010",
                      Input( 6) WHEN "00011",
                      Input( 7) WHEN "00100",
                      Input( 8) WHEN "00101",
                      Input( 9) WHEN "00110",
                      Input(10) WHEN "00111",
                      Input(11) WHEN "01000",
                      Input(12) WHEN "01001",
                      Input(13) WHEN "01010",
                      Input(14) WHEN "01011",
                      Input(15) WHEN "01100",
                      Input(16) WHEN "01101",
                      Input(17) WHEN "01110",
                      Input(18) WHEN "01111",
                      Input(19) WHEN "10000",
                      Input(20) WHEN "10001",
                      Input(21) WHEN "10010",
                      Input(22) WHEN "10011",
                      Input(23) WHEN "10100",
                      Input(24) WHEN "10101",
                      Input(25) WHEN "10110",
                      Input(26) WHEN "10111",
                      Input(27) WHEN "11000",
                      Input(28) WHEN "11001",
                      Input(29) WHEN "11010",
                      Input(30) WHEN "11011",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 4) <= Input( 4) WHEN "00000",
                      Input( 5) WHEN "00001",
                      Input( 6) WHEN "00010",
                      Input( 7) WHEN "00011",
                      Input( 8) WHEN "00100",
                      Input( 9) WHEN "00101",
                      Input(10) WHEN "00110",
                      Input(11) WHEN "00111",
                      Input(12) WHEN "01000",
                      Input(13) WHEN "01001",
                      Input(14) WHEN "01010",
                      Input(15) WHEN "01011",
                      Input(16) WHEN "01100",
                      Input(17) WHEN "01101",
                      Input(18) WHEN "01110",
                      Input(19) WHEN "01111",
                      Input(20) WHEN "10000",
                      Input(21) WHEN "10001",
                      Input(22) WHEN "10010",
                      Input(23) WHEN "10011",
                      Input(24) WHEN "10100",
                      Input(25) WHEN "10101",
                      Input(26) WHEN "10110",
                      Input(27) WHEN "10111",
                      Input(28) WHEN "11000",
                      Input(29) WHEN "11001",
                      Input(30) WHEN "11010",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 5) <= Input( 5) WHEN "00000",
                      Input( 6) WHEN "00001",
                      Input( 7) WHEN "00010",
                      Input( 8) WHEN "00011",
                      Input( 9) WHEN "00100",
                      Input(10) WHEN "00101",
                      Input(11) WHEN "00110",
                      Input(12) WHEN "00111",
                      Input(13) WHEN "01000",
                      Input(14) WHEN "01001",
                      Input(15) WHEN "01010",
                      Input(16) WHEN "01011",
                      Input(17) WHEN "01100",
                      Input(18) WHEN "01101",
                      Input(19) WHEN "01110",
                      Input(20) WHEN "01111",
                      Input(21) WHEN "10000",
                      Input(22) WHEN "10001",
                      Input(23) WHEN "10010",
                      Input(24) WHEN "10011",
                      Input(25) WHEN "10100",
                      Input(26) WHEN "10101",
                      Input(27) WHEN "10110",
                      Input(28) WHEN "10111",
                      Input(29) WHEN "11000",
                      Input(30) WHEN "11001",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 6) <= Input( 6) WHEN "00000",
                      Input( 7) WHEN "00001",
                      Input( 8) WHEN "00010",
                      Input( 9) WHEN "00011",
                      Input(10) WHEN "00100",
                      Input(11) WHEN "00101",
                      Input(12) WHEN "00110",
                      Input(13) WHEN "00111",
                      Input(14) WHEN "01000",
                      Input(15) WHEN "01001",
                      Input(16) WHEN "01010",
                      Input(17) WHEN "01011",
                      Input(18) WHEN "01100",
                      Input(19) WHEN "01101",
                      Input(20) WHEN "01110",
                      Input(21) WHEN "01111",
                      Input(22) WHEN "10000",
                      Input(23) WHEN "10001",
                      Input(24) WHEN "10010",
                      Input(25) WHEN "10011",
                      Input(26) WHEN "10100",
                      Input(27) WHEN "10101",
                      Input(28) WHEN "10110",
                      Input(29) WHEN "10111",
                      Input(30) WHEN "11000",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 7) <= Input( 7) WHEN "00000",
                      Input( 8) WHEN "00001",
                      Input( 9) WHEN "00010",
                      Input(10) WHEN "00011",
                      Input(11) WHEN "00100",
                      Input(12) WHEN "00101",
                      Input(13) WHEN "00110",
                      Input(14) WHEN "00111",
                      Input(15) WHEN "01000",
                      Input(16) WHEN "01001",
                      Input(17) WHEN "01010",
                      Input(18) WHEN "01011",
                      Input(19) WHEN "01100",
                      Input(20) WHEN "01101",
                      Input(21) WHEN "01110",
                      Input(22) WHEN "01111",
                      Input(23) WHEN "10000",
                      Input(24) WHEN "10001",
                      Input(25) WHEN "10010",
                      Input(26) WHEN "10011",
                      Input(27) WHEN "10100",
                      Input(28) WHEN "10101",
                      Input(29) WHEN "10110",
                      Input(30) WHEN "10111",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 8) <= Input( 8) WHEN "00000",
                      Input( 9) WHEN "00001",
                      Input(10) WHEN "00010",
                      Input(11) WHEN "00011",
                      Input(12) WHEN "00100",
                      Input(13) WHEN "00101",
                      Input(14) WHEN "00110",
                      Input(15) WHEN "00111",
                      Input(16) WHEN "01000",
                      Input(17) WHEN "01001",
                      Input(18) WHEN "01010",
                      Input(19) WHEN "01011",
                      Input(20) WHEN "01100",
                      Input(21) WHEN "01101",
                      Input(22) WHEN "01110",
                      Input(23) WHEN "01111",
                      Input(24) WHEN "10000",
                      Input(25) WHEN "10001",
                      Input(26) WHEN "10010",
                      Input(27) WHEN "10011",
                      Input(28) WHEN "10100",
                      Input(29) WHEN "10101",
                      Input(30) WHEN "10110",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith( 9) <= Input( 9) WHEN "00000",
                      Input(10) WHEN "00001",
                      Input(11) WHEN "00010",
                      Input(12) WHEN "00011",
                      Input(13) WHEN "00100",
                      Input(14) WHEN "00101",
                      Input(15) WHEN "00110",
                      Input(16) WHEN "00111",
                      Input(17) WHEN "01000",
                      Input(18) WHEN "01001",
                      Input(19) WHEN "01010",
                      Input(20) WHEN "01011",
                      Input(21) WHEN "01100",
                      Input(22) WHEN "01101",
                      Input(23) WHEN "01110",
                      Input(24) WHEN "01111",
                      Input(25) WHEN "10000",
                      Input(26) WHEN "10001",
                      Input(27) WHEN "10010",
                      Input(28) WHEN "10011",
                      Input(29) WHEN "10100",
                      Input(30) WHEN "10101",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(10) <= Input(10) WHEN "00000",
                      Input(11) WHEN "00001",
                      Input(12) WHEN "00010",
                      Input(13) WHEN "00011",
                      Input(14) WHEN "00100",
                      Input(15) WHEN "00101",
                      Input(16) WHEN "00110",
                      Input(17) WHEN "00111",
                      Input(18) WHEN "01000",
                      Input(19) WHEN "01001",
                      Input(20) WHEN "01010",
                      Input(21) WHEN "01011",
                      Input(22) WHEN "01100",
                      Input(23) WHEN "01101",
                      Input(24) WHEN "01110",
                      Input(25) WHEN "01111",
                      Input(26) WHEN "10000",
                      Input(27) WHEN "10001",
                      Input(28) WHEN "10010",
                      Input(29) WHEN "10011",
                      Input(30) WHEN "10100",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(11) <= Input(11) WHEN "00000",
                      Input(12) WHEN "00001",
                      Input(13) WHEN "00010",
                      Input(14) WHEN "00011",
                      Input(15) WHEN "00100",
                      Input(16) WHEN "00101",
                      Input(17) WHEN "00110",
                      Input(18) WHEN "00111",
                      Input(19) WHEN "01000",
                      Input(20) WHEN "01001",
                      Input(21) WHEN "01010",
                      Input(22) WHEN "01011",
                      Input(23) WHEN "01100",
                      Input(24) WHEN "01101",
                      Input(25) WHEN "01110",
                      Input(26) WHEN "01111",
                      Input(27) WHEN "10000",
                      Input(28) WHEN "10001",
                      Input(29) WHEN "10010",
                      Input(30) WHEN "10011",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(12) <= Input(12) WHEN "00000",
                      Input(13) WHEN "00001",
                      Input(14) WHEN "00010",
                      Input(15) WHEN "00011",
                      Input(16) WHEN "00100",
                      Input(17) WHEN "00101",
                      Input(18) WHEN "00110",
                      Input(19) WHEN "00111",
                      Input(20) WHEN "01000",
                      Input(21) WHEN "01001",
                      Input(22) WHEN "01010",
                      Input(23) WHEN "01011",
                      Input(24) WHEN "01100",
                      Input(25) WHEN "01101",
                      Input(26) WHEN "01110",
                      Input(27) WHEN "01111",
                      Input(28) WHEN "10000",
                      Input(29) WHEN "10001",
                      Input(30) WHEN "10010",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(13) <= Input(13) WHEN "00000",
                      Input(14) WHEN "00001",
                      Input(15) WHEN "00010",
                      Input(16) WHEN "00011",
                      Input(17) WHEN "00100",
                      Input(18) WHEN "00101",
                      Input(19) WHEN "00110",
                      Input(20) WHEN "00111",
                      Input(21) WHEN "01000",
                      Input(22) WHEN "01001",
                      Input(23) WHEN "01010",
                      Input(24) WHEN "01011",
                      Input(25) WHEN "01100",
                      Input(26) WHEN "01101",
                      Input(27) WHEN "01110",
                      Input(28) WHEN "01111",
                      Input(29) WHEN "10000",
                      Input(30) WHEN "10001",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(14) <= Input(14) WHEN "00000",
                      Input(15) WHEN "00001",
                      Input(16) WHEN "00010",
                      Input(17) WHEN "00011",
                      Input(18) WHEN "00100",
                      Input(19) WHEN "00101",
                      Input(20) WHEN "00110",
                      Input(21) WHEN "00111",
                      Input(22) WHEN "01000",
                      Input(23) WHEN "01001",
                      Input(24) WHEN "01010",
                      Input(25) WHEN "01011",
                      Input(26) WHEN "01100",
                      Input(27) WHEN "01101",
                      Input(28) WHEN "01110",
                      Input(29) WHEN "01111",
                      Input(30) WHEN "10000",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(15) <= Input(15) WHEN "00000",
                      Input(16) WHEN "00001",
                      Input(17) WHEN "00010",
                      Input(18) WHEN "00011",
                      Input(19) WHEN "00100",
                      Input(20) WHEN "00101",
                      Input(21) WHEN "00110",
                      Input(22) WHEN "00111",
                      Input(23) WHEN "01000",
                      Input(24) WHEN "01001",
                      Input(25) WHEN "01010",
                      Input(26) WHEN "01011",
                      Input(27) WHEN "01100",
                      Input(28) WHEN "01101",
                      Input(29) WHEN "01110",
                      Input(30) WHEN "01111",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(16) <= Input(16) WHEN "00000",
                      Input(17) WHEN "00001",
                      Input(18) WHEN "00010",
                      Input(19) WHEN "00011",
                      Input(20) WHEN "00100",
                      Input(21) WHEN "00101",
                      Input(22) WHEN "00110",
                      Input(23) WHEN "00111",
                      Input(24) WHEN "01000",
                      Input(25) WHEN "01001",
                      Input(26) WHEN "01010",
                      Input(27) WHEN "01011",
                      Input(28) WHEN "01100",
                      Input(29) WHEN "01101",
                      Input(30) WHEN "01110",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(17) <= Input(17) WHEN "00000",
                      Input(18) WHEN "00001",
                      Input(19) WHEN "00010",
                      Input(20) WHEN "00011",
                      Input(21) WHEN "00100",
                      Input(22) WHEN "00101",
                      Input(23) WHEN "00110",
                      Input(24) WHEN "00111",
                      Input(25) WHEN "01000",
                      Input(26) WHEN "01001",
                      Input(27) WHEN "01010",
                      Input(28) WHEN "01011",
                      Input(29) WHEN "01100",
                      Input(30) WHEN "01101",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(18) <= Input(18) WHEN "00000",
                      Input(19) WHEN "00001",
                      Input(20) WHEN "00010",
                      Input(21) WHEN "00011",
                      Input(22) WHEN "00100",
                      Input(23) WHEN "00101",
                      Input(24) WHEN "00110",
                      Input(25) WHEN "00111",
                      Input(26) WHEN "01000",
                      Input(27) WHEN "01001",
                      Input(28) WHEN "01010",
                      Input(29) WHEN "01011",
                      Input(30) WHEN "01100",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(19) <= Input(19) WHEN "00000",
                      Input(20) WHEN "00001",
                      Input(21) WHEN "00010",
                      Input(22) WHEN "00011",
                      Input(23) WHEN "00100",
                      Input(24) WHEN "00101",
                      Input(25) WHEN "00110",
                      Input(26) WHEN "00111",
                      Input(27) WHEN "01000",
                      Input(28) WHEN "01001",
                      Input(29) WHEN "01010",
                      Input(30) WHEN "01011",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(20) <= Input(20) WHEN "00000",
                      Input(21) WHEN "00001",
                      Input(22) WHEN "00010",
                      Input(23) WHEN "00011",
                      Input(24) WHEN "00100",
                      Input(25) WHEN "00101",
                      Input(26) WHEN "00110",
                      Input(27) WHEN "00111",
                      Input(28) WHEN "01000",
                      Input(29) WHEN "01001",
                      Input(30) WHEN "01010",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(21) <= Input(21) WHEN "00000",
                      Input(22) WHEN "00001",
                      Input(23) WHEN "00010",
                      Input(24) WHEN "00011",
                      Input(25) WHEN "00100",
                      Input(26) WHEN "00101",
                      Input(27) WHEN "00110",
                      Input(28) WHEN "00111",
                      Input(29) WHEN "01000",
                      Input(30) WHEN "01001",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(22) <= Input(22) WHEN "00000",
                      Input(23) WHEN "00001",
                      Input(24) WHEN "00010",
                      Input(25) WHEN "00011",
                      Input(26) WHEN "00100",
                      Input(27) WHEN "00101",
                      Input(28) WHEN "00110",
                      Input(29) WHEN "00111",
                      Input(30) WHEN "01000",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(23) <= Input(23) WHEN "00000",
                      Input(24) WHEN "00001",
                      Input(25) WHEN "00010",
                      Input(26) WHEN "00011",
                      Input(27) WHEN "00100",
                      Input(28) WHEN "00101",
                      Input(29) WHEN "00110",
                      Input(30) WHEN "00111",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(24) <= Input(24) WHEN "00000",
                      Input(25) WHEN "00001",
                      Input(26) WHEN "00010",
                      Input(27) WHEN "00011",
                      Input(28) WHEN "00100",
                      Input(29) WHEN "00101",
                      Input(30) WHEN "00110",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(25) <= Input(25) WHEN "00000",
                      Input(26) WHEN "00001",
                      Input(27) WHEN "00010",
                      Input(28) WHEN "00011",
                      Input(29) WHEN "00100",
                      Input(30) WHEN "00101",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(26) <= Input(26) WHEN "00000",
                      Input(27) WHEN "00001",
                      Input(28) WHEN "00010",
                      Input(29) WHEN "00011",
                      Input(30) WHEN "00100",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(27) <= Input(27) WHEN "00000",
                      Input(28) WHEN "00001",
                      Input(29) WHEN "00010",
                      Input(30) WHEN "00011",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(28) <= Input(28) WHEN "00000",
                      Input(29) WHEN "00001",
                      Input(30) WHEN "00010",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(29) <= Input(29) WHEN "00000",
                      Input(30) WHEN "00001",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(30) <= Input(30) WHEN "00000",
                      Input(31) WHEN OTHERS ;

WITH Shamt SELECT
ShiftRghtArith(31) <= Input(31) WHEN OTHERS ;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

END MainArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.Shifter(MainArch)
--PORT MAP   (Input    => SLV,
--            Shamt    => SLV,
--            ArithRlN => SLV,
--            Output   => SLV
--           );
------------------------------------------------------------------------------------------