------------------------------------------------------------------------------------------
--                                                                                      --
--                              Ivan Ricardo Diaz Gamarra                               --
--                                                                                      --
--  Project:                                                                            --
--  Date:                                                                               --
--                                                                                      --
------------------------------------------------------------------------------------------
--                                                                                      --
--                                                                                      --
--                                                                                      --
--                                                                                      --
------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BasicPackage.ALL;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ENTITY MainMemoryTestbench IS
    
    PORT   (DataRd     : IN  uint32;
            Address    : IN  uint32;
            RdWrEnable : IN  uint02;
            DataWr     : OUT uint32 
           );
    
END ENTITY MainMemoryTestbench;

------------------------------------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------------------------------------

ARCHITECTURE TbArch OF MainMemoryTestbench IS

SIGNAL Tmp : uint32;

BEGIN

------------------------------------------------------------
-- 
-- 
-- 
------------------------------------------------------------

WITH RdWrEnable SELECT
DataWr <= Tmp         WHEN "10",
          Tmp         WHEN "11",
          x"FFFFFFFF" WHEN OTHERS;

WITH Address SELECT
Tmp    <= "00001011000000000000010101101111" WHEN (Int2Slv(000,32)),
          "00001011000000000000010101101111" WHEN (Int2Slv(000,32)),
          "10000000000000000000111000110111" WHEN (Int2Slv(016,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(017,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(018,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(019,32)),
          "11111111101011100001111011110011" WHEN (Int2Slv(020,32)),
          "00000000001000000000010101101111" WHEN (Int2Slv(021,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(022,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(023,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(024,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(025,32)),
          "00011101000000000000000001100111" WHEN (Int2Slv(026,32)),
          "00000000000000000000000010110111" WHEN (Int2Slv(032,32)),
          "00000000000000000000111110110111" WHEN (Int2Slv(033,32)),
          "01111000011110000000011110110111" WHEN (Int2Slv(034,32)),
          "00011100000000000000000001100111" WHEN (Int2Slv(035,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(036,32)),
          "11111111101100001001010111110011" WHEN (Int2Slv(048,32)),
          "00010000000000000001101010110111" WHEN (Int2Slv(049,32)),
          "00010000000000000001101100110111" WHEN (Int2Slv(050,32)),
          "00010000000000000001101110110111" WHEN (Int2Slv(051,32)),
          "00010000000000000001110000110111" WHEN (Int2Slv(052,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(053,32)),
          "00100000000000000010101010110111" WHEN (Int2Slv(064,32)),
          "00100000000000000010101100110111" WHEN (Int2Slv(065,32)),
          "00100000000000000010101110110111" WHEN (Int2Slv(066,32)),
          "00100000000000000010110000110111" WHEN (Int2Slv(067,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(068,32)),
          "00110000000000000011101010110111" WHEN (Int2Slv(080,32)),
          "00110000000000000011101100110111" WHEN (Int2Slv(081,32)),
          "00110000000000000011101110110111" WHEN (Int2Slv(082,32)),
          "00110000000000000011110000110111" WHEN (Int2Slv(083,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(084,32)),
          "01000000000000000100101010110111" WHEN (Int2Slv(096,32)),
          "01000000000000000100101100110111" WHEN (Int2Slv(097,32)),
          "01000000000000000100101110110111" WHEN (Int2Slv(098,32)),
          "01000000000000000100110000110111" WHEN (Int2Slv(099,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(100,32)),
          "00010000000100000001101010110111" WHEN (Int2Slv(112,32)),
          "00010000000100000001101100110111" WHEN (Int2Slv(113,32)),
          "00010000000100000001101110110111" WHEN (Int2Slv(114,32)),
          "00010000000100000001110000110111" WHEN (Int2Slv(115,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(116,32)),
          "00100000000100000010101010110111" WHEN (Int2Slv(128,32)),
          "00100000000100000010101100110111" WHEN (Int2Slv(129,32)),
          "00100000000100000010101110110111" WHEN (Int2Slv(130,32)),
          "00100000000100000010110000110111" WHEN (Int2Slv(131,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(132,32)),
          "00110000000100000011101010110111" WHEN (Int2Slv(144,32)),
          "00110000000100000011101100110111" WHEN (Int2Slv(145,32)),
          "00110000000100000011101110110111" WHEN (Int2Slv(146,32)),
          "00110000000100000011110000110111" WHEN (Int2Slv(147,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(148,32)),
          "01000000000100000100101010110111" WHEN (Int2Slv(160,32)),
          "01000000000100000100101100110111" WHEN (Int2Slv(161,32)),
          "01000000000100000100101110110111" WHEN (Int2Slv(162,32)),
          "01000000000100000100110000110111" WHEN (Int2Slv(163,32)),
          "00110000001000000000000001110011" WHEN (Int2Slv(164,32)),
          "00000000000000000001010110110111" WHEN (Int2Slv(176,32)),
          "11111111111111111111011000110111" WHEN (Int2Slv(177,32)),
          "00000000000000011111011010110111" WHEN (Int2Slv(178,32)),
          "10101010101010101010011100110111" WHEN (Int2Slv(179,32)),
          "01010101010101010101011110110111" WHEN (Int2Slv(180,32)),
          "00000000000000010001100000110111" WHEN (Int2Slv(181,32)),
          "10000000000000000000100010110111" WHEN (Int2Slv(182,32)),
          "00000000110001011101000010010011" WHEN (Int2Slv(183,32)),
          "00000000110001100101000100010011" WHEN (Int2Slv(184,32)),
          "00000000000001100101111110010011" WHEN (Int2Slv(185,32)),
          "10101010101000000000100100110111" WHEN (Int2Slv(186,32)),
          "00000000110001101101000110010011" WHEN (Int2Slv(187,32)),
          "00000000110001110101001000010011" WHEN (Int2Slv(188,32)),
          "00000000110001111101001010010011" WHEN (Int2Slv(189,32)),
          "00000000110010000101001100010011" WHEN (Int2Slv(190,32)),
          "11111111111100000000111110010011" WHEN (Int2Slv(191,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(192,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(193,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(194,32)),
          "00000000010010010000001110110011" WHEN (Int2Slv(195,32)),
          "01000001000111111000111100110011" WHEN (Int2Slv(196,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(197,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(198,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(199,32)),
          "00000000000000000001010100010111" WHEN (Int2Slv(200,32)),
          "00001110000100000000010100010011" WHEN (Int2Slv(201,32)),
          "00000000000000001000010100010011" WHEN (Int2Slv(202,32)),
          "11111111111100001000010100010011" WHEN (Int2Slv(203,32)),
          "00000000000100000010010100010011" WHEN (Int2Slv(204,32)),
          "11111111111100000010010100010011" WHEN (Int2Slv(205,32)),
          "01111111111100000010010100010011" WHEN (Int2Slv(206,32)),
          "00000000000000000010010100010011" WHEN (Int2Slv(207,32)),
          "00000010000000011010010100010011" WHEN (Int2Slv(208,32)),
          "00000000000000001010010100010011" WHEN (Int2Slv(209,32)),
          "00000000000100000011010100010011" WHEN (Int2Slv(210,32)),
          "11111111111100000011010100010011" WHEN (Int2Slv(211,32)),
          "01111111111100000011010100010011" WHEN (Int2Slv(212,32)),
          "00000000000000000011010100010011" WHEN (Int2Slv(213,32)),
          "00000010000000011011010100010011" WHEN (Int2Slv(214,32)),
          "00000000000000001011010100010011" WHEN (Int2Slv(215,32)),
          "00000000001100001100010100010011" WHEN (Int2Slv(216,32)),
          "00000000001100001110010100010011" WHEN (Int2Slv(217,32)),
          "00000000001100001111010100010011" WHEN (Int2Slv(218,32)),
          "00000000001100001001010100010011" WHEN (Int2Slv(219,32)),
          "00000000000011111101010100010011" WHEN (Int2Slv(220,32)),
          "00000000000111111101010100010011" WHEN (Int2Slv(221,32)),
          "00000000100011111101010100010011" WHEN (Int2Slv(222,32)),
          "00000001111111111101010100010011" WHEN (Int2Slv(223,32)),
          "01000000000000111101010100010011" WHEN (Int2Slv(224,32)),
          "01000000000100111101010100010011" WHEN (Int2Slv(225,32)),
          "01000000100000111101010100010011" WHEN (Int2Slv(226,32)),
          "01000001111100111101010100010011" WHEN (Int2Slv(227,32)),
          "00000000010100100000010100110011" WHEN (Int2Slv(228,32)),
          "01000000000100000000010110110011" WHEN (Int2Slv(229,32)),
          "01000000101100000000010110110011" WHEN (Int2Slv(230,32)),
          "01000000000000000000010110110011" WHEN (Int2Slv(231,32)),
          "01000000011000011000010110110011" WHEN (Int2Slv(232,32)),
          "00000000000100001001010100110011" WHEN (Int2Slv(233,32)),
          "00000000011000001001010100110011" WHEN (Int2Slv(234,32)),
          "00000000001100001001010100110011" WHEN (Int2Slv(235,32)),
          "00000001111100001001010100110011" WHEN (Int2Slv(236,32)),
          "00000001111100000010010100110011" WHEN (Int2Slv(237,32)),
          "00000000000100000010010100110011" WHEN (Int2Slv(238,32)),
          "00000000001100110010010100110011" WHEN (Int2Slv(239,32)),
          "00000001111000110010010100110011" WHEN (Int2Slv(240,32)),
          "00000000000000001010010100110011" WHEN (Int2Slv(241,32)),
          "00000001111100000011010100110011" WHEN (Int2Slv(242,32)),
          "00000000000100000011010100110011" WHEN (Int2Slv(243,32)),
          "00000000001100110011010100110011" WHEN (Int2Slv(244,32)),
          "00000001111000110011010100110011" WHEN (Int2Slv(245,32)),
          "00000000000000001011010100110011" WHEN (Int2Slv(246,32)),
          "00000000001000100100010110110011" WHEN (Int2Slv(247,32)),
          "00000000010000100100010110110011" WHEN (Int2Slv(248,32)),
          "00000000001000100110010110110011" WHEN (Int2Slv(249,32)),
          "00000000010000100110010110110011" WHEN (Int2Slv(250,32)),
          "00000000001000100111010110110011" WHEN (Int2Slv(251,32)),
          "00000000010000100111010110110011" WHEN (Int2Slv(252,32)),
          "00000000000111111101010100110011" WHEN (Int2Slv(253,32)),
          "00000000011011111101010100110011" WHEN (Int2Slv(254,32)),
          "00000000001111111101010100110011" WHEN (Int2Slv(255,32)),
          "00000001111111111101010100110011" WHEN (Int2Slv(256,32)),
          "01000000000111111101010100110011" WHEN (Int2Slv(257,32)),
          "01000000011011111101010100110011" WHEN (Int2Slv(258,32)),
          "01000001111111111101010100110011" WHEN (Int2Slv(259,32)),
          "01000000000111111101010100110011" WHEN (Int2Slv(260,32)),
          "00000010000000001000011000110011" WHEN (Int2Slv(261,32)),
          "00000011111100001000011000110011" WHEN (Int2Slv(262,32)),
          "00000010001100110000011000110011" WHEN (Int2Slv(263,32)),
          "00000011111111111000011000110011" WHEN (Int2Slv(264,32)),
          "00000011111011111000011000110011" WHEN (Int2Slv(265,32)),
          "00000011111111110000011000110011" WHEN (Int2Slv(266,32)),
          "00000011111011110000011000110011" WHEN (Int2Slv(267,32)),
          "00000010000000001001011010110011" WHEN (Int2Slv(268,32)),
          "00000011111100001001011010110011" WHEN (Int2Slv(269,32)),
          "00000010001100110001011010110011" WHEN (Int2Slv(270,32)),
          "00000011111111111001011010110011" WHEN (Int2Slv(271,32)),
          "00000011111011111001011010110011" WHEN (Int2Slv(272,32)),
          "00000011111111110001011010110011" WHEN (Int2Slv(273,32)),
          "00000011111011110001011010110011" WHEN (Int2Slv(274,32)),
          "00000010000000001010011010110011" WHEN (Int2Slv(275,32)),
          "00000011111100001010011010110011" WHEN (Int2Slv(276,32)),
          "00000010001100110010011010110011" WHEN (Int2Slv(277,32)),
          "00000011111111111010011010110011" WHEN (Int2Slv(278,32)),
          "00000011111011111010011010110011" WHEN (Int2Slv(279,32)),
          "00000011111111110010011010110011" WHEN (Int2Slv(280,32)),
          "00000011111011110010011010110011" WHEN (Int2Slv(281,32)),
          "00000010000000001011011010110011" WHEN (Int2Slv(282,32)),
          "00000011111100001011011010110011" WHEN (Int2Slv(283,32)),
          "00000010001100110011011010110011" WHEN (Int2Slv(284,32)),
          "00000011111111111011011010110011" WHEN (Int2Slv(285,32)),
          "00000011111011111011011010110011" WHEN (Int2Slv(286,32)),
          "00000011111111110011011010110011" WHEN (Int2Slv(287,32)),
          "00000011111011110011011010110011" WHEN (Int2Slv(288,32)),
          "00000010000000001100011010110011" WHEN (Int2Slv(289,32)),
          "00000010000000001101011000110011" WHEN (Int2Slv(290,32)),
          "00000010000000001110010110110011" WHEN (Int2Slv(291,32)),
          "00000010000000001111011010110011" WHEN (Int2Slv(292,32)),
          "00000000000100001001010100010011" WHEN (Int2Slv(293,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(294,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(295,32)),
          "00000000000100001001010110010011" WHEN (Int2Slv(296,32)),
          "00000000000101011001010110010011" WHEN (Int2Slv(297,32)),
          "00000000000101011001010110010011" WHEN (Int2Slv(298,32)),
          "00000000000101011001010110010011" WHEN (Int2Slv(299,32)),
          "00000000000100001001011000010011" WHEN (Int2Slv(300,32)),
          "00000000000101100001011000010011" WHEN (Int2Slv(301,32)),
          "00000000000101100001011000010011" WHEN (Int2Slv(302,32)),
          "00000000000101100001011000010011" WHEN (Int2Slv(303,32)),
          "00000000000101100001011000010011" WHEN (Int2Slv(304,32)),
          "00000000000100001001010100010011" WHEN (Int2Slv(305,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(306,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(307,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(308,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(309,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(310,32)),
          "00110000000100101001010111110011" WHEN (Int2Slv(311,32)),
          "00110000010000101001010111110011" WHEN (Int2Slv(312,32)),
          "00110000010100001001010111110011" WHEN (Int2Slv(313,32)),
          "00110100001000101001010111110011" WHEN (Int2Slv(314,32)),
          "00110100001100101001010111110011" WHEN (Int2Slv(315,32)),
          "11110001001000101001010111110011" WHEN (Int2Slv(316,32)),
          "11110001001100101001010111110011" WHEN (Int2Slv(317,32)),
          "11110001010000101001010111110011" WHEN (Int2Slv(318,32)),
          "11111111101000101001010111110011" WHEN (Int2Slv(319,32)),
          "11111111101100101001010111110011" WHEN (Int2Slv(320,32)),
          "11111111110000101001010111110011" WHEN (Int2Slv(321,32)),
          "11111111110011111010011001110011" WHEN (Int2Slv(322,32)),
          "11111111110011111011011001110011" WHEN (Int2Slv(323,32)),
          "11111111110000000010011001110011" WHEN (Int2Slv(324,32)),
          "11111111110011111010011001110011" WHEN (Int2Slv(325,32)),
          "11111111110000000011011001110011" WHEN (Int2Slv(326,32)),
          "11111111101100000101011011110011" WHEN (Int2Slv(327,32)),
          "11111111110000000110011011110011" WHEN (Int2Slv(328,32)),
          "11111111101100000111011011110011" WHEN (Int2Slv(329,32)),
          "11111111110000000110011011110011" WHEN (Int2Slv(330,32)),
          "11111111101100000110011011110011" WHEN (Int2Slv(331,32)),
          "11111111110100000111011011110011" WHEN (Int2Slv(332,32)),
          "00011100011100000000100000100011" WHEN (Int2Slv(333,32)),
          "00011100011100000001100010100011" WHEN (Int2Slv(334,32)),
          "00011100011100000010100100100011" WHEN (Int2Slv(335,32)),
          "00000000011000000000010100000011" WHEN (Int2Slv(336,32)),
          "00000000011100000000010100000011" WHEN (Int2Slv(337,32)),
          "00000000100000000000010100000011" WHEN (Int2Slv(338,32)),
          "00000000011000000001010100000011" WHEN (Int2Slv(339,32)),
          "00000000011100000001010100000011" WHEN (Int2Slv(340,32)),
          "00000000100000000001010100000011" WHEN (Int2Slv(341,32)),
          "00000000011000000010010100000011" WHEN (Int2Slv(342,32)),
          "00000000011100000010010100000011" WHEN (Int2Slv(343,32)),
          "00000000100000000010010100000011" WHEN (Int2Slv(344,32)),
          "00000000011000000100010100000011" WHEN (Int2Slv(345,32)),
          "00000000011100000100010100000011" WHEN (Int2Slv(346,32)),
          "00000000100000000100010100000011" WHEN (Int2Slv(347,32)),
          "00000000011000000101010100000011" WHEN (Int2Slv(348,32)),
          "00000000011100000101010100000011" WHEN (Int2Slv(349,32)),
          "00000000100000000101010100000011" WHEN (Int2Slv(350,32)),
          "00000110000100000000000011100011" WHEN (Int2Slv(351,32)),
          "00000110001100011001000001100011" WHEN (Int2Slv(352,32)),
          "00000100011000011100111111100011" WHEN (Int2Slv(353,32)),
          "00000100001100110101111101100011" WHEN (Int2Slv(354,32)),
          "00000100001111111110111011100011" WHEN (Int2Slv(355,32)),
          "00000101111100011111111001100011" WHEN (Int2Slv(356,32)),
          "00000000000000000000010111100011" WHEN (Int2Slv(357,32)),
          "00010110011000000000000001100111" WHEN (Int2Slv(358,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(368,32)),
          "00010111000100000000000001100111" WHEN (Int2Slv(369,32)),
          "00000000000000000000111101100011" WHEN (Int2Slv(370,32)),
          "00010111001100000000000001100111" WHEN (Int2Slv(371,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(372,32)),
          "00010111010100000000000001100111" WHEN (Int2Slv(373,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(374,32)),
          "00010111011100000000000001100111" WHEN (Int2Slv(375,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(376,32)),
          "00010111100100000000000001100111" WHEN (Int2Slv(377,32)),
          "00000000000000000000001101100011" WHEN (Int2Slv(378,32)),
          "00010111101100000000000001100111" WHEN (Int2Slv(379,32)),
          "00000000000000001000000101100011" WHEN (Int2Slv(384,32)),
          "00000000000000000000111111100011" WHEN (Int2Slv(385,32)),
          "00011000001000000000000001100111" WHEN (Int2Slv(386,32)),
          "00000000000000001000001001100011" WHEN (Int2Slv(387,32)),
          "00000000000000001000000111100011" WHEN (Int2Slv(388,32)),
          "00000000000000001000000101100011" WHEN (Int2Slv(389,32)),
          "00000000000000000000111101100011" WHEN (Int2Slv(390,32)),
          "00011000011100000000000001100111" WHEN (Int2Slv(391,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(400,32)),
          "00011001000100000000000001100111" WHEN (Int2Slv(401,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(402,32)),
          "00011001001000000000000001100111" WHEN (Int2Slv(403,32)),
          "11111110000000000000000001100011" WHEN (Int2Slv(404,32)),
          "00011001010100000000000001100111" WHEN (Int2Slv(405,32)),
          "00000000000000001000000111100011" WHEN (Int2Slv(416,32)),
          "00000000000000001000000101100011" WHEN (Int2Slv(417,32)),
          "11111110000000000000000011100011" WHEN (Int2Slv(418,32)),
          "00011010001100000000000001100111" WHEN (Int2Slv(419,32)),
          "00000000000000001000001011100011" WHEN (Int2Slv(420,32)),
          "00000000000000001000001001100011" WHEN (Int2Slv(421,32)),
          "00000000000000001000000111100011" WHEN (Int2Slv(422,32)),
          "00000000000000001000000101100011" WHEN (Int2Slv(423,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(424,32)),
          "00011010100100000000000001100111" WHEN (Int2Slv(425,32)),
          "00000000000000001000001011100011" WHEN (Int2Slv(426,32)),
          "00000000000000001000001001100011" WHEN (Int2Slv(427,32)),
          "00000000000000001000000111100011" WHEN (Int2Slv(428,32)),
          "00000000000000001000000101100011" WHEN (Int2Slv(429,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(430,32)),
          "00011010111100000000000001100111" WHEN (Int2Slv(431,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(432,32)),
          "00011011000100000000000001100111" WHEN (Int2Slv(433,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(434,32)),
          "00110000010011111001011011110011" WHEN (Int2Slv(435,32)),
          "00000000000000000000011001100011" WHEN (Int2Slv(436,32)),
          "00011100000000000000000001100111" WHEN (Int2Slv(448,32)),
          "00000000000000000001010110110111" WHEN (Int2Slv(464,32)),
          "11111111111111111111011000110111" WHEN (Int2Slv(465,32)),
          "00000000000000011111011010110111" WHEN (Int2Slv(466,32)),
          "10101010101010101010011100110111" WHEN (Int2Slv(467,32)),
          "01010101010101010101011110110111" WHEN (Int2Slv(468,32)),
          "00000000000000010001100000110111" WHEN (Int2Slv(469,32)),
          "10000000000000000000100010110111" WHEN (Int2Slv(470,32)),
          "00000000110001011101000010010011" WHEN (Int2Slv(471,32)),
          "00000000110001100101000100010011" WHEN (Int2Slv(472,32)),
          "00000000000001100101111110010011" WHEN (Int2Slv(473,32)),
          "10101010101000000000100100110111" WHEN (Int2Slv(474,32)),
          "00000000110001101101000110010011" WHEN (Int2Slv(475,32)),
          "00000000110001110101001000010011" WHEN (Int2Slv(476,32)),
          "00000000110001111101001010010011" WHEN (Int2Slv(477,32)),
          "00000000110010000101001100010011" WHEN (Int2Slv(478,32)),
          "11111111111100000000111110010011" WHEN (Int2Slv(479,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(480,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(481,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(482,32)),
          "00000000010010010000001110110011" WHEN (Int2Slv(483,32)),
          "01000001000111111000111100110011" WHEN (Int2Slv(484,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(485,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(486,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(487,32)),
          "00001110000100000000010100010011" WHEN (Int2Slv(488,32)),
          "00000000000000001000010100010011" WHEN (Int2Slv(489,32)),
          "00000000000000001011010100110011" WHEN (Int2Slv(490,32)),
          "00000000001000100100010110110011" WHEN (Int2Slv(491,32)),
          "00000000000100001001010110010011" WHEN (Int2Slv(492,32)),
          "00000000000101010001010100010011" WHEN (Int2Slv(493,32)),
          "00000001111100011111000101100011" WHEN (Int2Slv(494,32)),
          "00000000000000000000000101100011" WHEN (Int2Slv(495,32)),
          "00011100000000000000000001100111" WHEN (Int2Slv(496,32)),
          "11111111101011100001111011110011" WHEN (Int2Slv(497,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(498,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(499,32)),
          "00000000000000000000000000110011" WHEN (Int2Slv(500,32)),
          "00001110000100000000010100010011" WHEN (Int2Slv(501,32)),
          "00000000000000001000010100010011" WHEN (Int2Slv(502,32)),
          "00011100000000000000000001100111" WHEN (Int2Slv(503,32)),
          "11111111111111111111111111111111" WHEN OTHERS;
END TbArch;

------------------------------------------------------------------------------------------
-- 
-- Summon This Block:
-- 
------------------------------------------------------------------------------------------
--BlockN: ENTITY WORK.MainMemoryTestbench(TbArch)
--PORT MAP   (DataRd     => SLV,
--            Address    => SLV,
--            RdWrEnable => SLV,
--            DataWr     => SLV
--           );
------------------------------------------------------------------------------------------
